module Decoder7Segment(
    input [3:0] in,
    output reg [6:0] seg
);
    always @(in) begin
        case(in)

        4'b0000: seg=7'b0000001; // active low logic display 0 on segment
        4'b0001: seg=7'b1001111; // 1
        4'b0010: seg=7'b0010010; // 2
        4'b0011: seg=7'b0000110; // 3
        4'b0100: seg=7'b1001100; // 4
        4'b0101: seg=7'b0100100; // 5
        4'b0110: seg=7'b0100000; // 6
        4'b0111: seg=7'b0001111; // 7
        4'b1000: seg=7'b0000000; // 8
        4'b1001: seg=7'b0001100; // 9
        endcase
    end


endmodule