module SevenSegDrive (
    input clk,
    input clr,
    input trigger,
    input [3:0] in1,
    input [3:0] in2,
    input [3:0] in3,
    input [3:0] in4,
    output reg [6:0] seg,
    output reg [3:0] an
);



endmodule